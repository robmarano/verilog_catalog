///////////////////////////////////////////////////////////////////////////////
//
// 2:1 multiplexer module
//
// A 2:1 mux module for your Computer Architecture Elements Catalog
//
// module: mux_2to1
// hdl: Verilog
//
// author: Your Name <your.name@cooper.edu>
//
///////////////////////////////////////////////////////////////////////////////

`ifndef MUX_2TO1
`define MUX_2TO1

module mux_2to1(add your module parameters here);
   //
   // ---------------- PORT DEFINITIONS ----------------
   //
   // ADD YOUR MODULE INPUTS AND OUTPUTS HERE

   //
   // ---------------- MODULE DESIGN IMPLEMENTATION ----------------
   //


endmodule

`endif // MUX_2TO1