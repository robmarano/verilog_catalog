///////////////////////////////////////////////////////////////////////////////
//
// D Flip Flow (DFF) module
//
// A DFF module for your Computer Architecture Elements Catalog
//
// module: dff
// hdl: Verilog
//
// author: Your Name <your.name@cooper.edu>
//
///////////////////////////////////////////////////////////////////////////////

`ifndef DFF
`define DFF

module dff(add your module parameters here);
   //
   // ---------------- PORT DEFINITIONS ----------------
   //
   // ADD YOUR MODULE INPUTS AND OUTPUTS HERE

   //
   // ---------------- MODULE DESIGN IMPLEMENTATION ----------------
   //

endmodule

`endif // DFF