///////////////////////////////////////////////////////////////////////////////
//
// 4:1 multiplexer module
//
// A 4:1 mux module for your Computer Architecture Elements Catalog
//
// module: mux_4to1
// hdl: Verilog
//
// author: Your Name <your.name@cooper.edu>
//
///////////////////////////////////////////////////////////////////////////////

`ifndef MUX_4TO1
`define MUX_4TO1

module mux_4to1(add your module parameters here);
   //
   // ---------------- PORT DEFINITIONS ----------------
   //
   // ADD YOUR MODULE INPUTS AND OUTPUTS HERE

   //
   // ---------------- MODULE DESIGN IMPLEMENTATION ----------------
   //

endmodule

`endif // MUX_4TO1