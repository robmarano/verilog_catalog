///////////////////////////////////////////////////////////////////////////////
//
// Counter module
//
// A counter module for your Computer Architecture Elements Catalog
//
// module: counter
// hdl: Verilog
//
// author: Your Name <your.name@cooper.edu>
//
///////////////////////////////////////////////////////////////////////////////

`ifndef COUNTER
`define COUNTER

module counter(add your module parameters here);
   //
   // ---------------- PORT DEFINITIONS ----------------
   //
   // ADD YOUR MODULE INPUTS AND OUTPUTS HERE

   //
   // ---------------- MODULE DESIGN IMPLEMENTATION ----------------
   //

endmodule

`endif // COUNTER