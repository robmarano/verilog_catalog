///////////////////////////////////////////////////////////////////////////////
//
// Shift Logical Right module
//
// A shift logical right (slr) module for your Computer Architecture Elements Catalog
//
// module: slr
// hdl: Verilog
//
// author: Your Name <your.name@cooper.edu>
//
///////////////////////////////////////////////////////////////////////////////

`ifndef SLR
`define SLR

module slr(add your module parameters here);
   //
   // ---------------- PORT DEFINITIONS ----------------
   //
   // ADD YOUR MODULE INPUTS AND OUTPUTS HERE

   //
   // ---------------- MODULE DESIGN IMPLEMENTATION ----------------
   //

endmodule

`endif // SLR