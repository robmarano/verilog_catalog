///////////////////////////////////////////////////////////////////////////////
//
// Sign Extender module
//
// A sign extension module for your Computer Architecture Elements Catalog
//
// module: signext
// hdl: Verilog
//
// author: Your Name <your.name@cooper.edu>
//
///////////////////////////////////////////////////////////////////////////////

`ifndef SIGNEXT
`define SIGNEXT

module signext(add your module parameters here);
   //
   // ---------------- PORT DEFINITIONS ----------------
   //
   // ADD YOUR MODULE INPUTS AND OUTPUTS HERE

   //
   // ---------------- MODULE DESIGN IMPLEMENTATION ----------------
   //

endmodule

`endif // SIGNEXT