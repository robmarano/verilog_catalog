///////////////////////////////////////////////////////////////////////////////
//
// Clock module
//
// A clock module for your Computer Architecture Elements Catalog
//
// module: clock
// hdl: Verilog
//
// author: Your Name <your.name@cooper.edu>
//
///////////////////////////////////////////////////////////////////////////////

`ifndef CLOCK
`define CLOCK

module clock(add your module parameters here);
   //
   // ---------------- PORT DEFINITIONS ----------------
   //
   // ADD YOUR MODULE INPUTS AND OUTPUTS HERE

   //
   // ---------------- MODULE DESIGN IMPLEMENTATION ----------------
   //

endmodule

`endif // CLOCK